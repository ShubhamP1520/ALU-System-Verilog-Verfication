package alu_pkg;
  //`include "alu.v"
  `include "alu_transaction.sv"
  `include "alu_generator.sv"
  `include "driver.sv"
  `include "alu_reference_model.sv"
  `include "alu_monitor.sv"
  `include "alu_scoreboard.sv"
  `include "alu_environment.sv"
  `include "alu_test.sv"
  //`include "alu.v"
endpackage
